-- reset generator
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity icds1813 is
  port(
    port1 : in std_ulogic;
    port2 : in std_ulogic;
    port3 : in std_ulogic
    );
end entity;

architecture rtl of icds1813 is
begin
end architecture;
