
module icds1813(
input wire port1 = 0,
input wire port2 = 0,
input wire port3 = 0
);

endmodule