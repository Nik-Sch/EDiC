-- 7segment display
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ic5082_7340 is
  port (
    port1 : in std_ulogic;
    port2 : in std_ulogic;
    port3 : in std_ulogic;
    port4 : in std_ulogic;
    port5 : in std_ulogic;
    port6 : in std_ulogic;
    port7 : in std_ulogic;
    port8 : in std_ulogic
    );
end entity;

architecture rtl of ic5082_7340 is
begin
-- currently no logic
end architecture;
