module icBerg40(
input wire port1,
input wire port2,
input wire port3,
input wire port4,
input wire port5,
output wire port6,
input wire port7,
output wire port8,
input wire port9,
output wire port10,
input wire port11,
output wire port12,
input wire port13,
output wire port14,
input wire port15,
output wire port16,
input wire port17,
output wire port18,
input wire port19,
output wire port20,
input wire port21,
output wire port22,
input wire port23,
output wire port24,
input wire port25,
output wire port26,
input wire port27,
output wire port28,
input wire port29,
output wire port30,
input wire port31,
output wire port32,
input wire port33,
output wire port34,
input wire port35,
output wire port36,
input wire port37,
input wire port38,
input wire port39,
input wire port40
);

assign port6 = port5;
assign port8 = port7;

assign port10 = port9;
assign port12 = port11;
assign port14 = port13;
assign port16 = port15;
assign port18 = port17;

assign port20 = port19;
assign port22 = port21;
assign port24 = port23;
assign port26 = port25;
assign port28 = port27;

assign port30 = port29;
assign port32 = port31;
assign port34 = port33;
assign port36 = port35;

endmodule