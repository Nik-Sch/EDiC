module icBerg10(
input wire port1,
input wire port2,
input wire port3,
output wire port4,
input wire port5,
output wire port6,
input wire port7,
output wire port8,
input wire port9,
input wire port10
);

assign port4 = port3;
assign port6 = port5;
assign port8 = port7;
endmodule