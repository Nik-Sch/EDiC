module icBerg26(
input wire port1,
input wire port2,
input wire port3,
input wire port4,
input wire port5,
output wire port6,
input wire port7,
output wire port8,
input wire port9,
output wire port10,
input wire port11,
output wire port12,
input wire port13,
output wire port14,
input wire port15,
output wire port16,
input wire port17,
output wire port18,
input wire port19,
output wire port20,
input wire port21,
output wire port22,
input wire port23,
input wire port24,
input wire port25,
input wire port26
);

assign port6 = port5;
assign port8 = port7;

assign port10 = port9;
assign port12 = port11;
assign port14 = port13;
assign port16 = port15;
assign port18 = port17;

assign port20 = port19;
assign port22 = port21;
endmodule;