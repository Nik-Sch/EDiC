module board_top(
  input wire i_clk100,

  // fpga buttons/switches
  input wire i_btnStep,
  input wire i_swInstrNCycle,
  input wire i_swStepNRun,
  input wire i_swEnableBreakpoint,
  input wire i_btnReset, // active low

  // included IO at 0xfe00
  output wire [7:0] o_cathodes, // dot + gfedcba
  output wire [7:0] o_anodes,
  input wire [9:0] i_switches,

  // expansion connector
  output reg [7:0] o_ramAddress,
  inout wire [7:0] io_bus,
  output reg o_ioNCE,
  output reg o_ctrlMemRamNOE,
  output reg o_nreset,
  output reg o_ctrlMemRamNWE,
  output reg o_clk,

  // tri-color led
  output reg o_ld17_r,
  output reg o_ld17_g,
  output reg o_ld17_b,

  // fpga debug
  output wire [7:0] o_r0,
  output wire [7:0] o_r1,

  // for included uart
  input wire i_serialIn,
  output wire o_serialOut
);

wire [7:0] s_expansionBusIn;
reg [7:0] s_expansionBusOut;
wire s_expansionBusNOE;
wire s_expansionIoNCE;
wire [7:0] s_expansionIoAddress;
wire s_expansionIoNOE;
wire s_expansionIoNWE;


reg [15:0] r_breakpoint;
reg r_breakpointSet;

wire s_resetn;
assign s_resetn = i_btnReset;

wire s_oszClk;
wire s_clkRam;
wire s_clkEEPROM;

clk_wiz_5Mhz inst_clk5Mhz(
  .clk_in1(i_clk100),
  .clk5(s_oszClk),
  .clkRam(s_clkRam),
  .clkEEPROM(s_clkEEPROM)
);

reg [1:0] r_oszClkDiv = 0;
always @(posedge s_oszClk) begin
  r_oszClkDiv <= r_oszClkDiv + 1;
end

reg [1:0] r_clkRamDiv = 2;
always @(posedge s_clkRam) begin
  r_clkRamDiv <= r_clkRamDiv + 1;
end

reg [1:0] r_clkEEPROMDiv = 3;
always @(posedge s_clkEEPROM) begin
  r_clkEEPROMDiv <= r_clkEEPROMDiv + 1;
end

always @(negedge s_oszClk, negedge s_resetn) begin
  r_breakpointSet <= 1;
  if (~r_breakpointSet) begin
    r_breakpoint <= {6'h00, i_switches};
  end

  if (~s_resetn) begin
    r_breakpointSet <= 0;
    r_breakpoint <= 0;
  end
end

generated inst_generated(
  .i_clk100(i_clk100),

  .i_oszClk(r_oszClkDiv[1]),
  .i_asyncRamSpecialClock(r_clkRamDiv[1]),
  .i_asyncEEPROMSpecialClock(r_clkEEPROMDiv[1]),
  .i_resetn(s_resetn),

  // button controls
  // 1 is closed, 0 is open
  .i_btnStep(i_btnStep),
  .i_swInstrNCycle(i_swInstrNCycle),
  .i_swStepNRun(i_swStepNRun),
  .i_swEnableBreakpoint(i_swEnableBreakpoint),
  .i_btnReset(~i_btnReset), // btn should be 1 if pressed -> active high
  .i_breakpointAddress(r_breakpoint),

  // expansion card
  .i_bus(s_expansionBusOut),
  .o_bus(s_expansionBusIn),
  .i_busNOE(s_expansionBusNOE),

  .o_ioNCE(s_expansionIoNCE),
  .o_ioAddress(s_expansionIoAddress),
  .o_ioNOE(s_expansionIoNOE),
  .o_ioNWE(s_expansionIoNWE),

  // fpga specific ports
  .o_cathodes(o_cathodes),
  .o_anodes(o_anodes),
  .i_switches(i_switches[7:0]),
  .o_r0(o_r0),
  .o_r1(o_r1)
);

// expansion_uart uart(
//   .i_clk100(i_clk100),
//   .i_clkDesign(r_clkRamDiv[1]),
//   .i_resetn(s_resetn),

//   .i_bus(s_expansionBusIn),
//   .o_bus(s_expansionBusOut),
//   .o_busNOE(s_expansionBusNOE),

//   .i_ioNCE(s_expansionIoNCE),
//   .i_ioAddress(s_expansionIoAddress),
//   .i_ioNOE(s_expansionIoNOE),
//   .i_ioNWE(s_expansionIoNWE),

//   .i_serialIn(i_serialIn),
//   .o_serialOut(o_serialOut)
// );
reg [7:0] io_bus_reg_out;
reg [7:0] io_bus_reg_in;

assign io_bus = (s_expansionIoNCE | s_expansionIoNOE) ? io_bus_reg_out : 8'hzz;
// assign s_expansionBusOut = (s_expansionIoNCE | s_expansionIoNOE) ? 8'hff : io_bus_reg_in;

// wire external expansion:
always @(posedge i_clk100) begin
  o_ramAddress <= s_expansionIoAddress;
  io_bus_reg_out <= s_expansionBusIn;
  io_bus_reg_in <= io_bus;
  s_expansionBusOut <= (s_expansionIoNCE | s_expansionIoNOE) ? 8'hff : io_bus_reg_in;
  o_ioNCE <= s_expansionIoNCE;
  o_ctrlMemRamNOE <= s_expansionIoNOE;
  o_nreset <= s_resetn;
  o_ctrlMemRamNWE <= s_expansionIoNWE;
  o_clk <= ~r_oszClkDiv[1];
end

endmodule