.title KiCad schematic
.include "/home/niklas/dev/KiCad-Spice-Library/Models/uncategorized/Bordodynovs Electronics Lib/sub/timers.lib"
XU1 GND /clock/thr /clock/clock +5V Net-_C1-Pad1_ /clock/thr /clock/dis +5V LM555
R2 /clock/thr /clock/dis 1k
R1 +5V /clock/dis 1k
V1 +5V GND 5V
R3 /clock/clock GND 10Meg
C1 Net-_C1-Pad1_ GND 0.01u
C2 /clock/thr GND 0.1u
.tran 1u 10m 0 uic 
.end
