// reset generator
module icds1813(
input wire port1,
input wire port2,
input wire port3
);

endmodule