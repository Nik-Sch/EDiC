
module ic28C256(
input wire port1 = 0,
input wire port2 = 0,
input wire port3 = 0,
input wire port4 = 0,
input wire port5 = 0,
input wire port6 = 0,
input wire port7 = 0,
input wire port8 = 0,
input wire port9 = 0,
input wire port10 = 0,
input wire port11 = 0,
input wire port12 = 0,
input wire port13 = 0,
input wire port14 = 0,
input wire port15 = 0,
input wire port16 = 0,
input wire port17 = 0,
input wire port18 = 0,
input wire port19 = 0,
input wire port20 = 0,
input wire port21 = 0,
input wire port22 = 0,
input wire port23 = 0,
input wire port24 = 0,
input wire port25 = 0,
input wire port26 = 0,
input wire port27 = 0,
input wire port28 = 0
);

endmodule