// 7segment display
module ic5082_7340(
input wire port1,
input wire port2,
input wire port3,
input wire port4,
input wire port5,
input wire port6,
input wire port7,
input wire port8
);

// currently no logic

endmodule